LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY CLK_DIVIDER IS
	GENERIC (PRE_SCALER : INTEGER := 8;
				COUNTER_BITS : INTEGER := 32);
	PORT (CLK_IN : IN STD_LOGIC;
			RESET_IN : IN STD_LOGIC;
		   CLK_OUT : OUT STD_LOGIC);
END CLK_DIVIDER;

ARCHITECTURE DIVIDER_LOGIC OF CLK_DIVIDER IS
	SIGNAL COUNTER_REG : STD_LOGIC_VECTOR (COUNTER_BITS-1 DOWNTO 0) := (OTHERS => '0');
	SIGNAL SIGNAL_OUT : STD_LOGIC := '0';
BEGIN
	PROCESS(CLK_IN)
	BEGIN
		IF (RESET_IN = '1') THEN
			COUNTER_REG <= (OTHERS => '0');
			SIGNAL_OUT <= '0';
		ELSIF (CLK_IN'EVENT AND CLK_IN = '1') THEN
			COUNTER_REG <= COUNTER_REG + '1';
			IF (TO_INTEGER(UNSIGNED(COUNTER_REG)) = PRE_SCALER) THEN
				SIGNAL_OUT <= NOT SIGNAL_OUT;
				COUNTER_REG <= (0 => '1', OTHERS => '0');
			END IF;
		END IF;
	END PROCESS;
	CLK_OUT <= SIGNAL_OUT;
END DIVIDER_LOGIC;